

module ALU (
  input clk,
  input rst,

  input [15:0] AC,
  input []
);

endmodule